module allgate(
  input a,b,
  output y1
);

  assign y1 = a&b;

endmodule